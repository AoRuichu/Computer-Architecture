module foward_unit#(
     parameter integer DATA_W     = 64 
)(
        
        input  wire [4:0] IF_ID_Rs1,
        input  wire [4:0] IF_ID_Rs2,
        input  wire       EX_MEM_reg_write,
        input  wire [4:0] EX_MEM_Rd,
        input  wire       MEM_WB_reg_write,
        input  wire [4:0] MEM_WB_Rd

);


endmodule;